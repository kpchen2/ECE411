module wb_stage
import rv32i_types::*;
(
    input   logic           clk,
    input   logic           rst,
    
    input   mem_wb_reg_t    mem_wb_reg
);

    always_comb begin
        
    end

endmodule : wb_stage